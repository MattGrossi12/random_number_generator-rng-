//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:47:20 04/02/2026 
// Design Name: 
// Module Name:    rng_control_path
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module rng_control_path(
    input clk_cp_i,
    input rst_cp_i,
    input req_card_state_cp,

    output state_o
);

//States:
localparam IDLE = 0;
localparam SEND = 1;

reg next_state;

always@(posedge clk_cp_i or negedge rst_cp_i)
    begin
        if(!rst_cp_i)
            begin
                next_state <= IDLE;
            end
        else 
        if(req_card_state_cp)
            begin 
                next_state <= SEND;
            end
        else
            begin
                next_state <= IDLE;
            end
    end

assign state_o = next_state;

endmodule